module unified_controller #(
    parameter GRID_WIDTH_X = 4,
    parameter GRID_WIDTH_Z = 1,
    parameter GRID_WIDTH_U = 3,
    parameter ITERATION_COUNTER_WIDTH = 8,  // counts to 255 iterations
    parameter MAXIMUM_DELAY = 3,
    parameter NUM_CONTEXTS = 2,
    parameter CTRL_FIFO_WIDTH = 64,
    parameter NUM_FPGAS = 5,
    parameter ROUTER_DELAY_COUNTER = 18,
    parameter LOGICAL_QUBITS_PER_DIM = 2
) (
    clk,
    reset,

    input_data,
    input_valid,
    input_ready,

    output_data,
    output_valid,
    output_ready,

    input_ctrl_rx_data,
    input_ctrl_rx_valid,
    input_ctrl_rx_ready,

    output_ctrl_tx_data,
    output_ctrl_tx_valid,
    output_ctrl_tx_ready,

    busy_PE, 
    odd_clusters_PE,
    measurements,
    correction,
    global_stage,

    router_busy,
    border_continous,
    FPGA_ID,
    measurement_fusion,
    reset_all_edges
);

`include "../../parameters/parameters.sv"

`define MAX(a, b) (((a) > (b)) ? (a) : (b))

localparam X_BIT_WIDTH = $clog2(GRID_WIDTH_X);
localparam Z_BIT_WIDTH = $clog2(GRID_WIDTH_Z);
localparam U_BIT_WIDTH = $clog2(GRID_WIDTH_U);
localparam FPGA_BIT_WIDTH = $clog2(NUM_FPGAS);
localparam ADDRESS_WIDTH = X_BIT_WIDTH + Z_BIT_WIDTH + U_BIT_WIDTH + FPGA_BIT_WIDTH;

localparam BYTES_PER_ROUND = ((GRID_WIDTH_X * GRID_WIDTH_Z  + 7) >> 3);
localparam ALIGNED_PU_PER_ROUND = (BYTES_PER_ROUND << 3);

localparam PU_COUNT_PER_ROUND = GRID_WIDTH_X * GRID_WIDTH_Z;
localparam PHYSICAL_GRID_WIDTH_U = (GRID_WIDTH_U % NUM_CONTEXTS == 0) ? 
                                   (GRID_WIDTH_U / NUM_CONTEXTS) : 
                                   (GRID_WIDTH_U / NUM_CONTEXTS + 1);

localparam PU_COUNT = PU_COUNT_PER_ROUND * PHYSICAL_GRID_WIDTH_U;

localparam NS_ERROR_COUNT_PER_ROUND = (GRID_WIDTH_X-1) * GRID_WIDTH_Z;
localparam EW_ERROR_COUNT_PER_ROUND = (GRID_WIDTH_X-1) * GRID_WIDTH_Z + 1;
localparam UD_ERROR_COUNT_PER_ROUND = GRID_WIDTH_X * GRID_WIDTH_Z;
localparam CORRECTION_COUNT_PER_ROUND = NS_ERROR_COUNT_PER_ROUND + EW_ERROR_COUNT_PER_ROUND + UD_ERROR_COUNT_PER_ROUND;

localparam BORDER_TOP_MSB = PU_COUNT - 1;
localparam BORDER_TOP_LSB = PU_COUNT_PER_ROUND * (PHYSICAL_GRID_WIDTH_U- 1);
localparam BORDER_BOT_MSB = PU_COUNT_PER_ROUND - 1;
localparam BORDER_BOT_LSB = 0;

localparam CTRL_MSG_MSB = 47;


input clk;
input reset;
output reg [STAGE_WIDTH-1:0] global_stage;
reg [STAGE_WIDTH-1:0] global_stage_previous;
reg [STAGE_WIDTH-1:0] global_stage_d;
reg [STAGE_WIDTH-1:0] global_stage_saved;
input [PU_COUNT - 1 : 0]  odd_clusters_PE;
input [PU_COUNT - 1 : 0]  busy_PE;
output reg [ALIGNED_PU_PER_ROUND-1:0] measurements;
input [CORRECTION_COUNT_PER_ROUND-1:0] correction;

input [7 : 0] input_data;
input input_valid;
output reg input_ready;

output reg [7 : 0] output_data;
output reg output_valid;
input output_ready;

input [CTRL_FIFO_WIDTH-1:0] input_ctrl_rx_data;
input input_ctrl_rx_valid;
output reg input_ctrl_rx_ready;

output reg [CTRL_FIFO_WIDTH-1:0] output_ctrl_tx_data;
output reg output_ctrl_tx_valid;
input output_ctrl_tx_ready;

input router_busy;
output reg [1:0] border_continous;
input [7:0] FPGA_ID;
output reg measurement_fusion;
output reg reset_all_edges;

reg result_valid;
reg [ITERATION_COUNTER_WIDTH-1:0] iteration_counter;
reg [31:0] cycle_counter;
reg [31:0] lower_half_counter;

reg busy;
reg odd_clusters;
reg border_busy;
reg [CONTEXT_COUNTER_WIDTH-1:0] current_context;

always@(posedge clk) begin
    busy <= |busy_PE;
    odd_clusters <= |odd_clusters_PE;
    border_busy <= |(busy_PE[BORDER_TOP_MSB : BORDER_TOP_LSB]) || |(busy_PE[BORDER_BOT_MSB : BORDER_BOT_LSB]);
end

reg[$clog2(ROUTER_DELAY_COUNTER+1)-1 : 0] router_busy_reg;

always@(posedge clk) begin
    if (reset) begin
        router_busy_reg <= 0;
    end else begin
        if(global_stage == STAGE_MERGE) begin
            if(router_busy) begin
                router_busy_reg <= ROUTER_DELAY_COUNTER;
            end else if( router_busy_reg > 0) begin
                router_busy_reg <= router_busy_reg - 1;
            end
        end else begin
            router_busy_reg <= 0;
        end
    end
end

// global_stage_d delayed logic
always @(posedge clk) begin
    if (reset) begin
        global_stage_d <= STAGE_IDLE;
    end else begin
        global_stage_d <= global_stage;
    end
end

reg cycle_counter_on;
reg cycle_counter_reset;

always @(posedge clk) begin
    if (reset) begin
        cycle_counter <= 0;
    end else begin
        if(cycle_counter_reset) begin
            cycle_counter <= 1; // By setting counter to 1 in a given cycle, we can ensure that the cycle counter always display the current cycle count instead of cycles elapsed. 
        end else if(cycle_counter_on) begin
            cycle_counter <= cycle_counter + 1;
        end
    end
end

always @(posedge clk) begin
    if (reset) begin
        global_stage_previous <= STAGE_IDLE;
    end else begin
        global_stage_previous <= global_stage;
    end
end

always@(*) begin
    if(global_stage == STAGE_GROW || global_stage == STAGE_MERGE || global_stage == STAGE_PEELING || global_stage == STAGE_RESET_ROOTS) begin
        cycle_counter_on = 1;
    end else if(global_stage == STAGE_WRITE_TO_MEM) begin
        if(global_stage_saved == STAGE_GROW || global_stage_saved == STAGE_MERGE || global_stage_saved == STAGE_PEELING || global_stage_saved == STAGE_RESET_ROOTS) begin
            cycle_counter_on = 1;
        end else begin
            cycle_counter_on = 0;
        end
    end else begin
        cycle_counter_on = 0;
    end
end

always@(*) begin
    if(global_stage == STAGE_IDLE && input_ctrl_rx_valid && input_ctrl_rx_ready && input_ctrl_rx_data [CTRL_MSG_MSB : CTRL_MSG_MSB - 7] == MEASUREMENT_DATA_HEADER && input_ctrl_rx_data [0] == 1'b0) begin // The last 0 is to ensure only to set it in the first stage
        cycle_counter_reset = 1;
    end else begin
        cycle_counter_reset = 0;
    end
end

always @(posedge clk) begin
    if (reset) begin
        iteration_counter <= 0;
    end else begin
        if (global_stage == STAGE_MEASUREMENT_LOADING) begin
            iteration_counter <= 0;
        end else if (global_stage == STAGE_GROW && global_stage_previous != STAGE_GROW) begin
            iteration_counter <= iteration_counter + 1;
        end
    end
end

always@(*) begin
    // Laksheen
    // if(measurement_fusion_stage == 2'b10) begin
    if(measurement_fusion_stage == 2'b01) begin
        measurement_fusion = 1;
    end else begin
        measurement_fusion = 0;
    end
end

localparam DELAY_COUNTER_WIDTH = $clog2(MAXIMUM_DELAY + 2);
reg [DELAY_COUNTER_WIDTH-1:0] delay_counter;

reg [15:0] messages_per_round_of_measurement;
reg [15:0] measurement_rounds;

wire [CORRECTION_COUNT_PER_ROUND - 1 : 0] output_fifo_data;
reg output_fifo_valid;
wire output_fifo_ready;

wire [CORRECTION_COUNT_PER_ROUND - 1 : 0] output_fifo_data_d;
wire output_fifo_valid_d;
wire output_fifo_ready_d;

reg [NUM_CONTEXTS -1 : 0] unsynced_merge;
reg [NUM_CONTEXTS -1 : 0] odd_clusters_in_context;
localparam CONTEXT_COUNTER_WIDTH = $clog2(NUM_CONTEXTS + 1);

reg measurement_fusion_on;
reg [1:0] measurement_fusion_stage; // 0 : First block, 1 : Second block, 3 : Merged block

reg fusion_on;
always@(*) begin
    if (reset) begin
        fusion_on = 0;
    end else begin
        if(NUM_CONTEXTS > 1 && (measurement_fusion_on==0 || (measurement_fusion_on == 1'b1 && measurement_fusion_stage == 2'b10))) begin
            fusion_on = 1;
        end else begin
            fusion_on = 0;
        end
    end
end


reg growing_incomplete; //Todo : In an optimized version use this. For the current version I'm not using it.

reg multi_fpga_mode;

always @(posedge clk) begin
    if (reset) begin
        global_stage <= STAGE_IDLE;
        delay_counter <= 0;
        result_valid <= 0;
        growing_incomplete <= 0;
        multi_fpga_mode <= 0;
        border_continous <= 2'b0;
        measurement_fusion_on <= 0;
        measurement_fusion_stage <= 0;
    end else begin
        case (global_stage)
            STAGE_IDLE: begin // 0
                if (input_ctrl_rx_valid && input_ctrl_rx_ready) begin
                    if(input_ctrl_rx_data [CTRL_MSG_MSB : CTRL_MSG_MSB - 7] == START_DECODING_MSG) begin
                        global_stage <= STAGE_PARAMETERS_LOADING;
                        delay_counter <= 0;
                        result_valid <= 0;
                        multi_fpga_mode <= input_ctrl_rx_data [0];
                        measurement_fusion_on <= input_ctrl_rx_data [1];
                        current_context <= 0; 
                        if(input_ctrl_rx_data[0] == 1'b1) begin
                            if(FPGA_ID != 1) begin
                                border_continous[0] <= 1'b1;
                            end
                            if(FPGA_ID != NUM_FPGAS - 1) begin
                                border_continous[1] <= 1'b1;
                            end
                        end
                    end else if(input_ctrl_rx_data [CTRL_MSG_MSB : CTRL_MSG_MSB - 7] == MEASUREMENT_DATA_HEADER) begin
                        global_stage <= STAGE_MEASUREMENT_PREPARING;
                        measurement_fusion_stage <= input_ctrl_rx_data [0];
                        current_context <= input_ctrl_rx_data [0];
                        delay_counter <= 0;
                        result_valid <= 0;
                        measurement_rounds <= 0;
                    end else if(input_ctrl_rx_data [CTRL_MSG_MSB : CTRL_MSG_MSB - 7] == MOVE_TO_STAGE) begin
                        global_stage <= STAGE_GROW;
                        delay_counter <= 0;
                        result_valid <= 0;
                    end
                end
            end

            STAGE_PARAMETERS_LOADING: begin // 6
                global_stage <= STAGE_IDLE;
                messages_per_round_of_measurement <= 0;
                measurement_rounds <= 0;
            end

            STAGE_MEASUREMENT_PREPARING: begin // 7
                if (input_valid && input_ready) begin
                    measurements[ALIGNED_PU_PER_ROUND-1:ALIGNED_PU_PER_ROUND-8] <= input_data;
                    if(ALIGNED_PU_PER_ROUND > 8) begin
                        measurements[ALIGNED_PU_PER_ROUND-9:0] <= measurements[ALIGNED_PU_PER_ROUND-1:8];
                    end
                    messages_per_round_of_measurement <= messages_per_round_of_measurement + 1;
                    if((messages_per_round_of_measurement + 1)*8 >= PU_COUNT_PER_ROUND) begin
                        global_stage <= STAGE_MEASUREMENT_LOADING;
                        delay_counter <= 0;
                        messages_per_round_of_measurement <= 0;
                        measurement_rounds <= measurement_rounds + 1;
                    end else begin
                        messages_per_round_of_measurement <= messages_per_round_of_measurement + 1;
                    end
                end
                unsynced_merge <= 0;
                odd_clusters_in_context <= 0;
            end

            STAGE_MEASUREMENT_LOADING: begin
                // Currently this is single cycle as only from external buffer happens.
                // In future might need multiple
                if(measurement_rounds < PHYSICAL_GRID_WIDTH_U) begin
                    global_stage <= STAGE_MEASUREMENT_PREPARING;
                    delay_counter <= 0;
                    result_valid <= 0;
                end else begin
                    global_stage_saved <= STAGE_MEASUREMENT_LOADING;
                    if(multi_fpga_mode == 1'b0) begin
                        if(!fusion_on) begin
                            global_stage <= STAGE_GROW;
                        end else begin
                            global_stage <= STAGE_WRITE_TO_MEM;
                        end
                    end else begin
                        global_stage <= STAGE_IDLE;
                    end
                    measurement_rounds <= 0;
                    delay_counter <= 0;
                    result_valid <= 0;
                end
            end

            STAGE_GROW: begin //2
                if(!fusion_on) begin
                    global_stage <= STAGE_MERGE;
                end else begin
                    global_stage <= STAGE_WRITE_TO_MEM;
                end
                global_stage_saved <= STAGE_GROW;
                delay_counter <= 0;
                measurement_rounds <= 0;
                growing_incomplete <= 1;
            end

            STAGE_MERGE: begin //3
                if (delay_counter >= MAXIMUM_DELAY) begin
                    if(multi_fpga_mode == 1'b0) begin
                        if(!busy) begin
                            delay_counter <= 0;
                            if(NUM_CONTEXTS == 1) begin
                                if(|odd_clusters == 1'b0) begin // everybody is even
                                    global_stage <= STAGE_PEELING;
                                end else begin // somebody is odd
                                    global_stage <= STAGE_GROW;
                                end
                            end else if(measurement_fusion_on && (measurement_fusion_stage == 2'b00 || measurement_fusion_stage == 2'b01)) begin
                                if(|odd_clusters == 1'b0) begin // everybody is even
                                    global_stage <= STAGE_WRITE_TO_MEM;
                                end else begin // somebody is odd
                                    global_stage <= STAGE_GROW;
                                end
                            end else begin
                                global_stage <= STAGE_WRITE_TO_MEM;
                            end
                            global_stage_saved <= STAGE_MERGE;
                            if(fusion_on) begin
                                odd_clusters_in_context[current_context] <= odd_clusters;
                            end  
                        end
                        if(border_busy) begin
                            if(fusion_on) begin
                                unsynced_merge[current_context] <= 1'b1;
                            end
                        end
                    end else begin
                        if (input_ctrl_rx_valid && input_ctrl_rx_ready && input_ctrl_rx_data [CTRL_MSG_MSB : CTRL_MSG_MSB - 7] == MOVE_TO_STAGE) begin
                            if(input_ctrl_rx_data[0] == 1'b0) begin
                                global_stage <= STAGE_PEELING;
                            end else begin
                                global_stage <= STAGE_GROW;
                            end
                        end
                    end
                end else begin
                    delay_counter <= delay_counter + 1;
                    unsynced_merge[current_context] <= 1'b0;
                end

            end           

            STAGE_PEELING: begin //4
                global_stage <= (NUM_CONTEXTS == 1 ? STAGE_RESULT_VALID : STAGE_WRITE_TO_MEM);
                global_stage_saved <= STAGE_PEELING;
            end

            STAGE_RESULT_VALID: begin //5
                measurement_rounds <= measurement_rounds + 1;
                if(measurement_rounds >= PHYSICAL_GRID_WIDTH_U - 1) begin
                    global_stage_saved <= STAGE_RESULT_VALID;
                    if(NUM_CONTEXTS == 1) begin
                        global_stage <= STAGE_IDLE;
                    end else begin
                        global_stage <= STAGE_WRITE_TO_MEM;
                    end
                    measurement_rounds <= 0;
                end
                delay_counter <= 0;
                result_valid <= 1;
            end

            STAGE_RESET_ROOTS: begin //8
                global_stage <= STAGE_WRITE_TO_MEM;
                global_stage_saved <= STAGE_RESET_ROOTS;
            end

            STAGE_WRITE_TO_MEM: begin //1
                if(fusion_on) begin
                    if(current_context < NUM_CONTEXTS -1) begin
                        if(global_stage_saved == STAGE_MERGE) begin
                            // if(growing_incomplete == 1'b1) begin
                            //     global_stage <= STAGE_GROW;
                            // end else begin
                            //     global_stage <= STAGE_MERGE;
                            // end
                            global_stage <= STAGE_MERGE;
                        end else if(global_stage_saved == STAGE_MEASUREMENT_LOADING) begin
                            global_stage <= STAGE_MEASUREMENT_PREPARING;
                        end else if(global_stage_saved == STAGE_PEELING) begin
                            global_stage <= STAGE_PEELING;
                        end else if(global_stage_saved == STAGE_RESULT_VALID) begin
                            global_stage <= STAGE_RESULT_VALID;
                        end else if(global_stage_saved == STAGE_GROW) begin
                            global_stage <= STAGE_GROW;
                        end else if(global_stage_saved == STAGE_RESET_ROOTS) begin
                            global_stage <= STAGE_RESET_ROOTS;
                        end
                        current_context <= current_context + 1;
                    end else begin
                        current_context <= 0;
                        growing_incomplete <= 0;
                        if(global_stage_saved == STAGE_MERGE) begin
                            if(|unsynced_merge == 1'b0) begin // everybody is synced
                                if(|odd_clusters_in_context == 1'b0) begin // everybody is even
                                    global_stage <= STAGE_PEELING;
                                end else begin // somebody is odd
                                    global_stage <= STAGE_GROW;
                                end
                            end else begin
                                global_stage <= STAGE_MERGE;
                            end
                        end else if(global_stage_saved == STAGE_MEASUREMENT_LOADING) begin
                            global_stage <= STAGE_GROW;
                        end else if(global_stage_saved == STAGE_PEELING) begin
                            global_stage <= STAGE_RESULT_VALID;
                        end else if(global_stage_saved == STAGE_RESULT_VALID) begin
                            global_stage <= STAGE_IDLE;
                        end else if(global_stage_saved == STAGE_GROW) begin
                            global_stage <= STAGE_MERGE;
                        end else if(global_stage_saved == STAGE_RESET_ROOTS) begin
                            global_stage <= STAGE_MERGE;
                        end
                    end
                // end else begin
                    delay_counter <= 0;
                // end
                end else begin
                    if(measurement_fusion_stage == 2'b00) begin
                        if(global_stage_saved == STAGE_MERGE) begin
                            global_stage <= STAGE_IDLE;
                            lower_half_counter <= cycle_counter;
                            current_context <= current_context + 1;
                        end
                    end else if(measurement_fusion_stage == 2'b01) begin
                        if(global_stage_saved == STAGE_MERGE) begin
                            global_stage <= STAGE_RESET_ROOTS;
                            measurement_fusion_stage <= 2'b10;
                            current_context <= 0;
                        end
                    end
                end
            end
            
            default: begin
                global_stage <= STAGE_IDLE;
            end
        endcase
    end
end

always@(*) begin
    if(global_stage == STAGE_MEASUREMENT_LOADING) begin
        if(measurement_fusion_on && measurement_fusion_stage != 2'b0) begin
            reset_all_edges = 0;
        end else begin
            reset_all_edges = 1;
        end
    end else begin
        reset_all_edges = 0;
    end
end

always@(*) begin
    if (reset) begin
        input_ready = 0;
    end else begin 
        if(global_stage == STAGE_MEASUREMENT_PREPARING) begin
            input_ready = 1;
        end else begin
            input_ready = 0;
        end
    end
end

always@(*) begin
    if (reset) begin
        output_fifo_valid = 0;
    end else begin 
        if(global_stage_d == STAGE_RESULT_VALID) begin
            output_fifo_valid = 1;
        end else begin
            output_fifo_valid = 0;
        end
    end
end

assign output_fifo_data = correction;

always@(*) begin
    if (reset) begin
        input_ctrl_rx_ready = 0;
    end else begin 
        if(global_stage == STAGE_IDLE) begin
            input_ctrl_rx_ready = 1;
        end else if(global_stage == STAGE_MERGE) begin
            if(multi_fpga_mode && delay_counter >= MAXIMUM_DELAY) begin
                input_ctrl_rx_ready = 1;
            end else begin
                input_ctrl_rx_ready = 0;
            end
        end else begin
            input_ctrl_rx_ready = 0;
        end
    end
end

reg result_is_send;

always@(posedge clk) begin
    if (reset) begin
        result_is_send <= 0;
    end else begin
        if(global_stage == STAGE_RESULT_VALID && current_context == 0) begin
            result_is_send <= 1;
        end else if(global_stage == STAGE_IDLE) begin
            result_is_send <= 0;
        end
    end
end

always@(*) begin
    output_ctrl_tx_valid = 0;
    output_ctrl_tx_valid = 0;
    output_ctrl_tx_data = 64'h0;
    if(reset) begin
        output_ctrl_tx_valid = 0;
    end else begin
        if(multi_fpga_mode == 1'b0) begin
            if(global_stage == STAGE_RESULT_VALID && result_is_send == 0) begin
                output_ctrl_tx_valid = 1;
                if(measurement_fusion_on) begin
                    output_ctrl_tx_data [CTRL_MSG_MSB : CTRL_MSG_MSB - 7] = lower_half_counter[7:0];
                end else begin
                    output_ctrl_tx_data [CTRL_MSG_MSB : CTRL_MSG_MSB - 7] = iteration_counter;
                end
                output_ctrl_tx_data [CTRL_MSG_MSB - 8 : CTRL_MSG_MSB - 23] = cycle_counter;
            end
        end else begin
            if(global_stage == STAGE_MERGE && delay_counter >= MAXIMUM_DELAY) begin
                if(input_ctrl_rx_valid && input_ctrl_rx_ready && input_ctrl_rx_data [CTRL_MSG_MSB : CTRL_MSG_MSB - 7] == SEND_ODD_AND_BUSY) begin
                    output_ctrl_tx_valid = 1;
                    output_ctrl_tx_data [CTRL_MSG_MSB : CTRL_MSG_MSB - 7] = NODE_RESULT_MSG;
                    output_ctrl_tx_data [1] = odd_clusters;
                    if(busy || router_busy_reg > 0) begin
                        output_ctrl_tx_data [0] = 1;
                    end else begin
                        output_ctrl_tx_data [0] = 0;
                    end
                end
            end
        end
    end
end

// FIFO
fifo_wrapper #(
    .WIDTH(CORRECTION_COUNT_PER_ROUND),
    .DEPTH(128)
) output_fifo (
    .clk(clk),
    .reset(reset),
    .input_data(output_fifo_data),
    .input_valid(output_fifo_valid),
    .input_ready(output_fifo_ready),
    .output_data(output_fifo_data_d),
    .output_valid(output_fifo_valid_d),
    .output_ready(output_fifo_ready_d)
);

wire [7 : 0] output_data_d2;
wire output_valid_d2;
reg output_ready_d2;

serializer #(
    .HUB_FIFO_WIDTH(CORRECTION_COUNT_PER_ROUND),
    .HUB_FIFO_PHYSICAL_WIDTH(8)
) output_serializer (
    .clk(clk),
    .reset(reset),
    .wide_fifo_data(output_fifo_data_d),
    .wide_fifo_valid(output_fifo_valid_d),
    .wide_fifo_ready(output_fifo_ready_d),
    .narrow_fifo_valid(output_valid_d2),
    .narrow_fifo_ready(output_ready_d2),
    .narrow_fifo_data(output_data_d2)
);

reg [31:0] output_message_counter;

always @(posedge clk) begin
    if (reset) begin
        output_message_counter <= 0;
    end else begin
        if(output_valid_d2 && output_ready) begin
            if(output_message_counter >= ((CORRECTION_COUNT_PER_ROUND + 7)>>3)*PHYSICAL_GRID_WIDTH_U*NUM_CONTEXTS + 2) begin
                output_message_counter <= 0;
            end else begin
                output_message_counter <= output_message_counter + 1;
            end
        end
    end
end

always@(*) begin
    case(output_message_counter)
        0: begin
            output_data = lower_half_counter[7:0];
            output_valid = output_valid_d2;
            output_ready_d2 = 0;
        end
        1: begin
            output_data = cycle_counter[15:8];
            output_valid = output_valid_d2;
            output_ready_d2 = 0;
        end
        2: begin
            output_data = cycle_counter[7:0];
            output_valid = output_valid_d2;
            output_ready_d2 = 0;
        end
        default: begin
            output_data = output_data_d2;
            output_valid = output_valid_d2;
            output_ready_d2 = output_ready;
        end
    endcase
end



endmodule